module And2bits(in0,in1,out);

output out;
input in0;
input in1;

assign out = in0&in1;

endmodule
